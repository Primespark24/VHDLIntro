------------------------------------------------
-- Module Name: majority4 
------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity majority4 is
-- complete the port statement for this module
end majority4;

architecture majority4 of majority4 is
begin
-- complete the behavioral code for this module
                             
end majority4;